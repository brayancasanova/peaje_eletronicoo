library verilog;
use verilog.vl_types.all;
entity Divisor_frecuencia is
    port(
        CLK             : in     vl_logic;
        out1            : out    vl_logic;
        out2            : out    vl_logic
    );
end Divisor_frecuencia;

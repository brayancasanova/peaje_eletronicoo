library verilog;
use verilog.vl_types.all;
entity peaje_eletronico_vlg_vec_tst is
end peaje_eletronico_vlg_vec_tst;

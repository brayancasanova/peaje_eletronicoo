library verilog;
use verilog.vl_types.all;
entity Divisor_frecuencia_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Divisor_frecuencia_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity Divisor_frecuencia_vlg_vec_tst is
end Divisor_frecuencia_vlg_vec_tst;

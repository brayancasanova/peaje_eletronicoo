library verilog;
use verilog.vl_types.all;
entity rom_5x5_vlg_vec_tst is
end rom_5x5_vlg_vec_tst;
